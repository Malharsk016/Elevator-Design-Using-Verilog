`timescale 1ns / 1ps

module elevatorproject_tf1;

    
      
endmodule
